package decrypt_pkg;
   import uvm_pkg::*;
`include "uvm_macros.svh"
   
   
`include "command_transaction.svh"   
`include "result_transaction.svh"
`include "coverage.svh"
`include "tester.svh"
`include "scoreboard.svh"
`include "driver.svh"
`include "command_monitor.svh"
`include "result_monitor.svh"
   
`include "env.svh"

`include "random_test.svh"
   
endpackage : decrypt_pkg
   